.title KiCad schematic
.include "setting/electronics/Simulation_SPICE.sp"
R8 Net-_C4-Pad1_ Net-_R8-Pad2_ 10kOhm
V6 0 Net-_U3-V-_ DC 15 
XU3 Net-_U3-+_ Net-_U3--_ Net-_U3-V+_ Net-_U3-V-_ Net-_R8-Pad2_ kicad_builtin_opamp POLE=300k GAIN=350 VOFF=0
R7 Net-_U3--_ Net-_C3-Pad1_ 100kOhm
R6 Net-_U3-+_ Net-_C3-Pad1_ 100kOhm
C4 Net-_C4-Pad1_ 0 100f
V5 Net-_U3-V+_ 0 DC 15 
R5 Net-_C4-Pad1_ 0 10kOhm
V8 Net-_C4-Pad1_ OUT4 TRNOISE( 10m 10p 0 0 0 0 0 ) AC 0 0 
C2 IN2 Net-_U1--_ 60f
R1 IN2 Net-_U1--_ 105kOhm
V2 0 Net-_U1-V-_ DC 15 
C6 IN2 Net-_U1--_ 68f
R3 Net-_U2--_ IN2 15kOhm
V1 Net-_U1-V+_ 0 DC 15 AC 1  
XU1 0 Net-_U1--_ Net-_U1-V+_ Net-_U1-V-_ IN2 kicad_builtin_opamp POLE=20Meg GAIN=1778 VOFF=0
C5 Net-_U3--_ IN3 100f
C3 Net-_C3-Pad1_ 0 100f
V4 0 Net-_U2-V-_ DC 15 
R4 IN3 Net-_U2--_ 150kOhm
V7 Net-_C3-Pad1_ 0 DC 1.5 AC 1  
V3 Net-_U2-V+_ 0 DC 15 
XU2 0 Net-_U2--_ Net-_U2-V+_ Net-_U2-V-_ IN3 kicad_builtin_opamp POLE=6.25Meg GAIN=251 VOFF=0
I1 0 IN1 PULSE( 0 0.3uA 0n 1p 1p 3.333n 1 0 ) AC 1  
C1 IN1 0 2.5p
R2 Net-_U1--_ IN1 1kOhm

.control
noise v(OUT4) V1 dec 100 100Hz 100GHz
* <output node> <source node *need to be with 'AC 1'*> 
* <point selection method> <number of points> 
* <frequency range start, need be with unit> <frequency range end> <noise generator contribution frequency>
setplot noise1
* plot with noise spectrum
wrdata output/afe/ABCStar_fe/noise.raw onoise_spectrum

tran 0.1n 100n
* <step> <stopping time>
wrdata output/afe/ABCStar_fe/tran.raw v(OUT4)
* save raw data
.endc

.end
