ucsc circuit 
* name of the circuit

* definition of BFR840L3RHESD, as a subcircuit
.subckt BFR840L3RHESD 1 2 3
*
Rcx 15 1 1.57895
Rbx 25 2 1.92983
Rex 35 3 0.0800447
*
CBEPAR 22 33 1.9449E-013
CBCPAR 22 11 3.44161E-014
CCEPAR 11 33 2.24848E-013
LB    22 20 3.04259E-010
LC   11 10  2.88058E-010
CBEPCK 20 30  1E-014
CBCPCK 20 10  1.5502E-014
CCEPCK 10 30  1E-014
LBX    20 25 9.04631E-011
LEX   30 35 3.71422E-011
LCX   10 15  9.15043E-011
*
R_CS_npn 55 5 500
*
D1 33 25 M_D1
D2 5 25  M_D2
*
R_NBL_fdb 22 25 3.2
R_PS 33 5 0.03
RSUB 30 5 0.03
*
D3 5 15 M_D3
D4 23 33 M_D4
D5 23 15 M_D5
*
R_NBL_e11g 15 11 1.8
*
Q1 11 22 33 55 M_BFR840L3RHESD
*
.MODEL M_D1 D(
+ IS=3E-015
+ N=1
+ RS=2.846
+ CJO=4E-014)
*
.MODEL M_D2 D(
+ IS=3E-015
+ N=1
+ RS=4170
+ CJO=4.5E-014)
*
.MODEL M_D3 D(
+ IS=6.911E-016
+ N=1.1
+ RS=1380
+ CJO =9.5E-014)
*
.MODEL M_D4 D(
+ IS=3.5E-015
+ N=1
+ RS=0.2
+ CJO =3E-014)
*
.MODEL M_D5 D(
+ IS=3.5E-015
+ N=1.02
+ RS=4.7
+ CJO =3E-014)
*
.MODEL 	M_BFR840L3RHESD	NPN(
+	TNOM = 25
+	IS	=	2.429E-016
+	BF	=	765.7
+	NF	=	1.012
+	VAF	=	375.1
+	IKF	=	0.0819
+	ISE	=	8.827E-014
+	NE	=	2.8
+	BR	=	194
+	NR	=	0.998
+	VAR	=	1.596
+	IKR	=	0.015
+	ISC	=	1.165E-015
+	NC	=	2
+	RB	=	7.53378
+	IRB	=	0
+	RBM	=	2.1
+	RE	=	0.4405
+	RC	=	7.246
+	XTB	=	-2.276
+	EG	=	1.11
+	XTI	=	-1.233
+	CJE	=	2.23E-014
+	VJE	=	0.9214
+	MJE	=	0.5
+	TF	=	1.1E-012
+	XTF	=	5.582
+	VTF	=	0.6828
+	ITF	=	0.4491
+	PTF	=	0.0214
+	CJC	=	6.6E-015
+	VJC	=	0.7723
+	MJC	=	1.005
+	XCJC	=	0.4894
+	TR	=	1E-010
+	CJS	=	1.147E-013
+	MJS	=	1.108
+   VJS =   0.6112
+	FC	=	0.578
+	KF	=	1.65E-011
+	AF	=	1.53)
.ends BFR840L3RHESD

I1 2 0 pulse(0 -10u 0 0.1n 1n 0.00000001n 20n 0)
* input current source
VCC 6 0 dc 2.25
* VCC, DC source
Rin 2 0 1MEG
* resistance of the sensor
C6 2 0 20p
* capacitance of the sensor
C1 2 3 3.3n
x1 5 3 0 BFR840L3RHESD
* the amplifier BFR840L3RHESD
R1 3 4 475
* feedback resistance
R2 4 5 3k
C2 4 5 3.3n
C5 5 out 3.3n
R4 out 0 50
L1 5 6 47U
R3 6 7 63.7
C7 8 0 10n
C8 7 0 10n
C3 7 0 1n
C4 7 0 1n
L2 8 7 2.2u
* some other devices

.control
tran 0.1p 20n
* <step> <stopping time>
wrdata ./raser/cflm/output/Current_test.raw v(out)
* save raw data
.endc

.end
